module day_2

fn test_level_1() {
	assert false
}

fn test_level_2() {
	assert false
}
