module day_3

fn test_level_1() {
	input := '467..114..
		...*......
		..35..633.
		......#...
		617*......
		.....+.58.
		..592.....
		......755.
		...$.*....
		+664.598.+
		.100...100'.replace('\t',
		'')

	solution := level_1(input)!
	assert solution == '4561'
}

fn test_level_2() {
	input := '467..114..
		...*......
		..35..633.
		......#...
		617*......
		.....+.58.
		..592.....
		......755.
		...$.*....
		+664.598.+'.replace('\t',
		'')

	solution := level_2(input)!
	assert solution == '467835'
}
