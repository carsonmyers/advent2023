module day_2

pub fn run(input string, level int) !string {
	if level == 1 {
		return level_1(input)
	} else {
		return level_2(input)
	}
}

fn level_1(input string) !string {
	return error('not implemented')
}

fn level_2(input string) !string {
	return error('not implemented')
}
