module day_5

fn test_level_1() {
	input := ''.replace('\t', '')

	solution := level_1(input)!
	assert solution == ''
}

fn test_level_2() {
	input := ''.replace('\t', '')

	solution := level_2(input)!
	assert solution == ''
}
