module main

// answer: POST https://adventofcode.com/:year/day/:day/answer { level: "1" | "2"; answer: string }